module Twos_comp #(parameter WIDTH = 6) (
    input  wire [WIDTH-1:0] data_in, 
    output wire [WIDTH-1:0] data_out  
);

    assign data_out = (~data_in) + 1'b1;

endmodule